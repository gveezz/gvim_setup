// Macro defines
`define

