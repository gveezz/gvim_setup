// $COMPONENT_NAME
// Headers include

module $COMPONENT_NAME # (
    // Configurable parameters
) (

);

// External functions and tasks
// Miscellaneous parameter task and functions

// Internal parameters (localparams)

// Registered outputs

// Virtually registered output (combinational regs)

// Internal registers

// Internal virtual registers (combinational regs)

// Internal wires

// Wires assignments

// Modules instantiations

// Testbench functionality

initial begin

   #0 ;
   
end

endmodule 
// end of $COMPONENT_NAME
