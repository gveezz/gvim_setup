////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////
//              Copyright $YEAR by KDPOF. All right reserved.
////////////////////////////////////////////////////////////////////////////////
// Component: $COMPONENT_NAME
// Date     : $Date: $
// Version  : $Revision: $
// Author   : SAZ
// Summary  : TODO: write summary
//            report bugs to simone.azzalin@kdpof.com 
////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////
// Macro defines
////////////////////////////////////////////////////////////////////////////////

`define 

// end of $COMPONENT_NAME
