// Macro defines
`define 

// end of $COMPONENT_NAME
