////////////////////////////////////////////////////////////////////////////////
// Headers include
////////////////////////////////////////////////////////////////////////////////

module $COMPONENT_NAME
(
   // System interface
   // -- inputs
   SClk,
   Reset_n,
   SyncRst,
   // Data interface
   // --inputs
   DataInVal,
   DataIn,
   // --outputs
   DataOutVal,
   DataOut
);

////////////////////////////////////////////////////////////////////////////////
// External functions and tasks
////////////////////////////////////////////////////////////////////////////////
// Miscellaneous parameter task and functions

////////////////////////////////////////////////////////////////////////////////
// Configurable parameters
////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////
// Internal parameters (localparams) that affect ports
////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////
// Module I/O
////////////////////////////////////////////////////////////////////////////////

input  logic SClk;       // COMMENT
input  logic Reset_n;    // COMMENT
input  logic SyncRst;    // COMMENT
input  logic DataInVal;  // COMMENT
input  logic DataIn;     // COMMENT
output logic DataOutVal; // COMMENT
output logic DataOut;    // COMMENT

////////////////////////////////////////////////////////////////////////////////
// Internal parameters (localparams)
////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////
// Registered outputs
////////////////////////////////////////////////////////////////////////////////

///////////////////////////////////////////////////////////////////////////////
// Virtually registered output (combinational regs)
////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////
// Internal registers
////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////
// Internal virtual registers (combinational regs)
////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////
// Internal wires
////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////
// Wires assignments
////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////
// Modules instantiations
////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////
// Module functionality
////////////////////////////////////////////////////////////////////////////////

always_comb begin

end

always_ff @(posedge SClk or negedge Reset_n) begin
   if (!Reset_n) begin
      DataOutVal <= 0;
      DataOut    <= 0;
   end else begin
      if (SyncRst) begin
         DataOutVal <= 0;
         DataOut    <= 0;
      end
   end
end

endmodule 
// end of $COMPONENT_NAME
