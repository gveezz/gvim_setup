`timescale 1ns/1ps
// Headers include

module $COMPONENT_NAME ();

// External functions and tasks
// Miscellaneous parameter task and functions

// Configurable parameters

// Internal parameters (localparams) that affect ports

// Module I/O

// Internal parameters (localparams)

// Registered outputs

// Virtually registered output (combinational regs)

// Internal registers

// Internal virtual registers (combinational regs)

// Internal wires

// Wires assignments

// Modules instantiations

// Testbench functionality

initial begin
   #0 ; 
end

endmodule 
// end of $COMPONENT_NAME
