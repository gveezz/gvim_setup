`timescale 1ns/1ps
// Headers include

module $COMPONENT_NAME # (
    // Configurable parameters
) ( 

);

// External functions and tasks

// Localparams

// Specparams

// Registered outputs

// Internal combinational regs

// Internal registers

// Internal wires

// Wires assignments

// Logic

// Real

// Modules instantiations

// Testbench functionality

initial begin
    #0 ; 
end

endmodule

