// Headers include

module $COMPONENT_NAME #(
   // Configurable parameters
   parameter DATA_W = 8
) (
   // System interface
   // -- inputs
   input logic SClk,
   input logic SyncRst,
   // Data interface
   // --inputs
   input logic DataInVal,
   input logic [DATA_W-1:0] DataIn,
   // --outputs
   output logic DataOutVal,
   output logic [DATA_W-1:0] DataOut
);

// External functions and tasks
// Miscellaneous parameter task and functions

// Configurable parameters

// Internal parameters (localparams)

// Module I/O

// Internal parameters (localparams)

// Registered outputs

// Virtually registered output (combinational regs)

// Internal registers

// Internal virtual registers (combinational regs)

// Internal wires

// Wires assignments

// Modules instantiations

// Module functionality

always_comb begin

end

always_ff @(posedge SClk) begin
   if (!SyncRst) begin
        DataOutVal <= 0;
        DataOut    <= 0;
   end else begin
        DataOutVal <= DataInVal;
        DataOut    <= DataIn;
   end
end

endmodule 

