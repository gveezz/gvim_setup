`timescale 1ns/1ps
// Headers include

module $COMPONENT_NAME # (
    // Configurable parameters
) (

);

// External functions and tasks
// Miscellaneous parameter task and functions

// Internal parameters (localparams)

// Registered outputs

// Virtually registered output (combinational regs)

// Internal registers

// Internal virtual registers (combinational regs)

// Internal wires

// Wires assignments

// Modules instantiations

// Testbench functionality

initial begin
    $dumpfile ("$COMPONENT_NAME.vcd");
    $dumpvars (0, $COMPONENT_NAME);
    #0 ;
end

endmodule 

