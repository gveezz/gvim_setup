// Macro defines
`define XXX

