////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////
//              Copyright 2024 by KDPOF. All right reserved.
////////////////////////////////////////////////////////////////////////////////
// Component: <Component name here>
// Date     : $Date: $
// Version  : $Revision: $
// Author   : SAZ
// Summary  : <Component summary here>
////////////////////////////////////////////////////////////////////////////////
////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////
// Headers include
////////////////////////////////////////////////////////////////////////////////

module module_name
(
   // System interface
   // -- inputs
   SClk,
   Reset_n,
   SyncRst,
   // Data interface
   // --inputs
   IDataVal,
   IData,
   // --outputs
   ODataVal,
   OData
);

////////////////////////////////////////////////////////////////////////////////
// External functions and tasks
////////////////////////////////////////////////////////////////////////////////
// Miscellaneous parameter task and functions

////////////////////////////////////////////////////////////////////////////////
// Configurable parameters
////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////
// Internal parameters (localparams) that affect ports
////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////
// Module I/O
////////////////////////////////////////////////////////////////////////////////

input  SClk;     // comment here
input  Reset_n;  // comment here
input  SyncRst;  // comment here
input  IDataVal; // comment here
input  IData;    // comment here
output ODataVal; // comment here
output OData;    // comment here

////////////////////////////////////////////////////////////////////////////////
// Internal parameters (localparams)
////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////
// Registered outputs
////////////////////////////////////////////////////////////////////////////////

reg ODataVal;
reg OData;

///////////////////////////////////////////////////////////////////////////////
// Virtually registered output (combinational regs)
////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////
// Internal registers
////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////
// Internal virtual registers (combinational regs)
////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////
// Internal wires
////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////
// Wires assignments
////////////////////////////////////////////////////////////////////////////////

////////////////////////////////////////////////////////////////////////////////
// Module description
////////////////////////////////////////////////////////////////////////////////

always @(posedge SClk or negedge Reset_n) begin
   if (!Reset_n) begin
      ODataVal <= 0;
      OData    <= 0;
   end else begin
      // handle sync clk logic here

      if (SyncRst) begin
         ODataVal <= 0;
         OData    <= 0;
      end
   end
end

endmodule

