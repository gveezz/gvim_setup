// $COMPONENT_NAME
// Macro defines
`define
// end of $COMPONENT_NAME
